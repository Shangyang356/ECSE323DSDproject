-- this circuit builds communications between three modules such as flash read control, altera up core, and audio interface.
-- 
-- entity name: g26_flash_read
--
-- Copyright (C) 2015 Chuan Qin, Wei Wang
-- Version 1.0
-- Author:  Chuan Qin; chuan.qin2@mail.mcgill.ca
--			Wei Wang; wei.wang18@mail.mcgill.ca
-- Date: March 16, 2015
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;



ENTITY g26_flash_read IS
GENERIC (
		FLASH_MEMORY_ADDRESS_WIDTH 	: INTEGER := 22;
		FLASH_MEMORY_DATA_WIDTH 		: INTEGER := 8
);
	PORT
	(	
		clk_50 			: IN std_logic; -- clk should be 50MHz 
		rst 			: IN std_logic;  
		shiftoctave     : in std_logic;
		volume			: in std_logic_vector (3 downto 0);
		trigger 		: IN std_logic; -- trigger = 1 resets the sample address to the beginning
		note			: IN unsigned(3 downto 0); -- selects the note to be played (within an octave)
		octave 			: IN unsigned(2 downto 0); -- the octave the note should be played at (4 octave range)
		sample_data 	: OUT std_logic_vector(15 downto 0); -- a single 16 bit sample value, to be sent to the audio codec chip
		--data_size_o 	: OUT unsigned(21 downto 0); -- number of samples in the wave file (for display on the LEDs)	
		
		i_data 			: IN STD_LOGIC_VECTOR(FLASH_MEMORY_DATA_WIDTH - 1 DOWNTO 0);			
		-- Signals to be connected to Flash chip via proper I/O ports
		FL_ADDR 		: OUT 	STD_LOGIC_VECTOR(FLASH_MEMORY_ADDRESS_WIDTH - 1 DOWNTO 0);
		FL_DQ 			: INOUT 	STD_LOGIC_VECTOR(FLASH_MEMORY_DATA_WIDTH - 1 DOWNTO 0);
		FL_CE_N,
		FL_OE_N,
		FL_WE_N,
		FL_RST_N 		: OUT 	STD_LOGIC;
		

		
		INIT 			: IN std_logic;
		AUD_MCLK 		: OUT std_logic; -- codec master clock input
		AUD_BCLK 		: OUT std_logic; -- digital audio bit clock
		AUD_DACDAT 		: OUT std_logic; -- DAC data lines
		AUD_DACLRCK 	: OUT std_logic; -- DAC data left/right select
		I2C_SDAT 		: OUT std_logic; -- serial interface data line
		I2C_SCLK 		: OUT std_logic  -- serial interface clock
	);
END g26_flash_read;

ARCHITECTURE func OF g26_flash_read IS

signal tempofo_data 			: std_logic_vector(7 downto 0);
signal tempofo_done 			: std_logic;
signal tempofflash_address 		: unsigned(21 downto 0);
signal tempofread_start 		: std_logic;
signal rippleouttemp1 			: std_logic;
signal rippleouttemp2 			: std_logic;
signal rippleouttemp3 			: std_logic;
signal rippleouttemp4 			: std_logic;
--signal tempofdata_size_o 		: unsigned (21 downto 0);
signal tempofpulse 				: std_logic;
signal tempofsample_data 		: std_logic_vector (15 downto 0);
signal temp1 					:std_logic_vector (23 downto 0);

component g26_flash_read_control
	port(
		clk_50 			: IN std_logic; -- clk should be 50MHz 
		rst 			: IN std_logic;  
		shiftoctave       : in std_logic;
		read_done 		: IN std_logic; -- indication from the flash memory that the read operation is complete
		step 			: IN std_logic;
		odata			: IN std_logic_vector(7 downto 0); -- output of the flash memory
		trigger 		: IN std_logic; -- trigger = 1 resets the sample address to the beginning
		note 			: IN unsigned(3 downto 0); -- selects the note to be played (within an octave)
		octave 			: IN unsigned(2 downto 0); -- the octave the note should be played at (4 octave range)
		flash_address 	: OUT unsigned(21 downto 0); -- address for the flash memory read operation
		read_start 		: OUT std_logic; -- request a read operation on the flash memory
		sample_data 	: OUT std_logic_vector(15 downto 0) -- a single 16 bit sample value, to be sent to the audio codec chip
		);
	end component;

component Altera_UP_Flash_Memory_UP_Core_Standalone
	port(
		i_clock 		: IN 		STD_LOGIC;
		i_reset_n 		: IN 		STD_LOGIC;
		i_address 		: IN 		STD_LOGIC_VECTOR(FLASH_MEMORY_ADDRESS_WIDTH - 1 DOWNTO 0);
		i_data 			: IN 		STD_LOGIC_VECTOR(FLASH_MEMORY_DATA_WIDTH - 1 DOWNTO 0);
		i_read,
		i_write,
		i_erase 		: IN 		STD_LOGIC;
		o_data 			: OUT 	STD_LOGIC_VECTOR(FLASH_MEMORY_DATA_WIDTH - 1 DOWNTO 0);
		o_done 			: OUT 	STD_LOGIC;
		
		-- Signals to be connected to Flash chip via proper I/O ports
		FL_ADDR 		: OUT 	STD_LOGIC_VECTOR(FLASH_MEMORY_ADDRESS_WIDTH - 1 DOWNTO 0);
		FL_DQ 			: INOUT 	STD_LOGIC_VECTOR(FLASH_MEMORY_DATA_WIDTH - 1 DOWNTO 0);
		FL_CE_N,
		FL_OE_N,
		FL_WE_N,
		FL_RST_N 		: OUT 	STD_LOGIC
		);
	end component;
	

component g26_audio_interface
	port(
		LDATA, RDATA	: IN signed(23 downto 0); -- parallel external data inputs
		clk 			: IN std_logic; -- clk should be 50MHz 
		rst 			: IN std_logic;  
		INIT			: IN std_logic;  
		W_EN			: IN std_logic;
		pulse 			: OUT std_logic; -- sample sync pulse
		AUD_MCLK 		: OUT std_logic; -- codec master clock input
		AUD_BCLK		: OUT std_logic; -- digital audio bit clock
		AUD_DACDAT      : OUT std_logic; -- DAC data lines
		AUD_DACLRCK 	: OUT std_logic; -- DAC data left/right select
		I2C_SDAT 		: OUT std_logic; -- serial interface data line
		I2C_SCLK 		: OUT std_logic  -- serial interface clock
	    );
	end component;

begin
	--data_size_o <= tempofdata_size_o;
	sample_data <= tempofsample_data;
	--temp1 <= std_LOGIC_VECTOR(TO_SIGNED(TO_INTEGER(signed(tempofsample_data)) *TO_INTEGER(unsigned(volume)),19)& "00000") ;
	temp1 <= tempofsample_data & "00000000";
	Gate1: g26_flash_read_control
	PORT MAP (
	clk_50 => clk_50,
	rst => not rst,
	shiftoctave => shiftoctave,
	read_done => tempofo_done,
	step => tempofpulse,
	odata => tempofo_data,
	trigger => not(trigger),
	note => note,
	octave => octave,
	flash_address => tempofflash_address,
	read_start => tempofread_start,
	sample_data => tempofsample_data
	);
	
	Gate2: Altera_UP_Flash_Memory_UP_Core_Standalone
	PORT MAP (
	i_clock => clk_50,
	i_reset_n => (rst),
	i_address => std_logic_vector(tempofflash_address),
	i_read => tempofread_start,
	i_data => i_data,
	i_write => '0',
	i_erase => '0',
	o_data => tempofo_data,
	o_done => tempofo_done,
	FL_ADDR => FL_ADDR,
	FL_DQ 	=> FL_DQ,
	FL_CE_N => FL_CE_N,
	FL_OE_N => FL_OE_N,
	FL_WE_N => FL_WE_N,
	FL_RST_N => FL_RST_N);
	
	
	Gate3: g26_audio_interface
	PORT MAP (
		clk => clk_50,
		rst => not rst,
		W_EN => '1',
		INIT => not INIT,
		LDATA => signed(temp1),
		RDATA => signed(temp1),
		pulse => tempofpulse,
		AUD_MCLK => AUD_MCLK,
		AUD_BCLK => AUD_BCLK,
		AUD_DACDAT => AUD_DACDAT,
		AUD_DACLRCK => AUD_DACLRCK,
		I2C_SDAT => I2C_SDAT,
		I2C_SCLK => I2C_SCLK
	);
end func;	
	